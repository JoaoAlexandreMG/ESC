module gnot16 (
    input [15:0] A,  
    output [15:0] Out  
);
    assign Out = ~A;
endmodule
