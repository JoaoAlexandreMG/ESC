module gor(
    input A, B,
    output Out
);
    assign Out = A | B;
endmodule
