module gxor(
    input A, B,
    output Y
);
    assign Y = A ^ B; 
endmodule